// Code your design here
module rom(
  output reg [3:0] data,
  input clk,
  input en,
  input [3:0] addr
);
  
  reg [3:0] rom[15:0];
  
  always@(posedge clk)
    begin
      if(en)
        data <= rom[addr];
      else
        data <= 4'bxxxx;
    end
  
  initial begin
      rom[0] = 4'b0010;
      rom[1] = 4'b0010;
      rom[2] = 4'b1110;
      rom[3] = 4'b0010;
      rom[4] = 4'b0100;
      rom[5] = 4'b1010;
      rom[6] = 4'b1100;
      rom[7] = 4'b0000;
      rom[8] = 4'b1010;
      rom[9] = 4'b0010;
      rom[10] = 4'b1110;
      rom[11] = 4'b0010;
      rom[12] = 4'b0100;
      rom[13] = 4'b1010;
      rom[14] = 4'b1100;
      rom[15] = 4'b0000;
  end
endmodule
